`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/11/09 15:33:32
// Design Name: 
// Module Name: des_E
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module des_E(
    input [31:0] R,
    output [47:0] expanded_R
    );

assign expanded_R = {
    R[31-31], R[31-0], R[31-1], R[31-2], R[31-3], R[31-4], 
    R[31-3], R[31-4], R[31-5], R[31-6], R[31-7], R[31-8],
    R[31-7], R[31-8], R[31-9], R[31-10], R[31-11], R[31-12],
    R[31-11], R[31-12], R[31-13], R[31-14], R[31-15], R[31-16],
    R[31-15], R[31-16], R[31-17], R[31-18], R[31-19], R[31-20],
    R[31-19], R[31-20], R[31-21], R[31-22], R[31-23], R[31-24],
    R[31-23], R[31-24], R[31-25], R[31-26], R[31-27], R[31-28],
    R[31-27], R[31-28], R[31-29], R[31-30], R[31-31], R[31-0]
};

endmodule
